ENTITY jurados IS
PORT ( 
