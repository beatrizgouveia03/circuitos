ENTITY reg IS
PORT (	d : IN BIT;
	clk : IN BIT;
	q : OUT BIT);
END reg;

